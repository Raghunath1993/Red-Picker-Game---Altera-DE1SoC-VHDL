library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;
use work.screen.all;
USE IEEE.math_real.all;

Entity sync is
PORT(
CLK: IN STD_LOGIC;
HSYNC,VSYNC:OUT STD_LOGIC;
R,G,B:OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
SWITCH: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
LED0: OUT STD_LOGIC
);
END sync;

ARCHITECTURE MAIN OF SYNC IS

SIGNAL HPOS: INTEGER RANGE 0 TO 800:=0;
SIGNAL VPOS: INTEGER RANGE 0 TO 525:=0;
--SIGNAL COLOR: INTEGER RANGE 0 TO 3:=0;
SIGNAL COUNTER16: INTEGER :=0;
SIGNAL LOCATION: STD_LOGIC_VECTOR(11 DOWNTO 0):= "100110101111"; 
SIGNAL RANDOM_NUMBER: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL REDPOS: STD_LOGIC_VECTOR(3 DOWNTO 0):="0111";
SIGNAL FLAG:STD_LOGIC:='0';
SIGNAL FFLAG:STD_LOGIC:='0';

COMPONENT RAND IS
PORT(
clk : in std_logic;
RANDOM_NUMBER : out std_logic_vector (3 downto 0));
END COMPONENT RAND;

BEGIN
C3: rand PORT MAP(clk,RANDOM_NUMBER);

PROCESS(CLK)
BEGIN
IF((SWITCH = REDPOS ) OR (SWITCH = "0001")) THEN
		FLAG <= '1';
		IF(COUNTER16 < 10) THEN
		   LED0 <= '0' ; 
			COUNTER16 <= COUNTER16 + 1;
			FFLAG <= '0';
		ELSE
		   LED0 <= '1' ;
		   FFLAG <= '1';
		END IF;
ELSE
		FLAG <='0';	
END IF;
		
	
IF(FLAG = '1') THEN
FLAG <= '0';
CASE RANDOM_NUMBER IS
WHEN "0000" => 
      LOCATION<="100110111101";
		REDPOS<="0111";
WHEN "0001" => 
      LOCATION<="100110101111";
		REDPOS<="0111";
WHEN "0010" => 
      LOCATION<="100111110101";
		REDPOS<="0111";
WHEN "0011" => 
      LOCATION<="100111101110";
		REDPOS<="0111";
WHEN "0100" => 
      LOCATION<="110100111101";
		REDPOS<="1011";
WHEN "0101" => 
      LOCATION<="110100101111";
		REDPOS<="1011";
WHEN "0110" => 
      LOCATION<="110101100111";
		REDPOS<="1101";
WHEN "0111" => 
      LOCATION<="110101111100";
		REDPOS<="1110";
WHEN "1000" => 
      LOCATION<="111100110101";
		REDPOS<="1011";
WHEN "1001" => 
      LOCATION<="111100101110";
		REDPOS<="1011";
WHEN "1010" => 
      LOCATION<="111110100101";
		REDPOS<="1101";
WHEN "1011" => 
      LOCATION<="111110101100";
		REDPOS<="1110";
WHEN "1100" => 
      LOCATION<="101100110111";
		REDPOS<="1011";
WHEN "1101" => 
      LOCATION<="101100111110";
		REDPOS<="1011";
WHEN "1110" => 
      LOCATION<="101110100111";
		REDPOS<="1101";
WHEN "1111" => 
      LOCATION<="101110111100";
		REDPOS<="1110";
END CASE;

END IF;
END PROCESS;



PROCESS(CLK)
--variable seed1,seed2: positive;
--variable rand: real;
--variable int_rand : integer;

BEGIN
  --uniform(seed1,seed2,rand);
  --int_rand := integer (rand*24);
  
  IF(CLK'EVENT AND CLK='1') THEN
	  IF (FFLAG ='0') THEN
			IF((HPOS>110 AND HPOS<210) AND(VPOS>70 AND VPOS<170)) THEN
				R<=(OTHERS=>LOCATION(11));
				G<=(OTHERS=>LOCATION(10));
				B<=(OTHERS=>LOCATION(9));
			ELSIF((HPOS>110 AND HPOS<210) AND(VPOS>310 AND VPOS<410)) THEN
				R<=(OTHERS=>LOCATION(8));
				G<=(OTHERS=>LOCATION(7));
				B<=(OTHERS=>LOCATION(6));
			ELSIF((HPOS>430 AND HPOS<530) AND(VPOS >70 AND VPOS<170)) THEN
				R<=(OTHERS=>LOCATION(5));
				G<=(OTHERS=>LOCATION(4));
				B<=(OTHERS=>LOCATION(3));
			ELSIF((HPOS>430 AND HPOS<530) AND(VPOS >310 AND VPOS<410)) THEN
				R<=(OTHERS=>LOCATION(2));
				G<=(OTHERS=>LOCATION(1));
				B<=(OTHERS=>LOCATION(0));
			ELSE
				R<=(OTHERS=>'0');
				G<=(OTHERS=>'0');
				B<=(OTHERS=>'0');
			END IF;
		ELSE
			IF((VPOS>70 AND VPOS<240) AND(HPOS>295 AND HPOS<345)) THEN
				R<=(OTHERS=>'1');
				G<=(OTHERS=>'0');
				B<=(OTHERS=>'0');
			ELSIF((HPOS>295 AND HPOS<345) AND(VPOS>260 AND VPOS<310)) THEN
				R<=(OTHERS=>'1');
				G<=(OTHERS=>'0');
				B<=(OTHERS=>'0');
			ELSE
				R<=(OTHERS=>'0');
				G<=(OTHERS=>'0');
				B<=(OTHERS=>'0');
			END IF;
	  END IF;
	
	IF(HPOS<800) THEN
		HPOS<=HPOS+1;
	ELSIF(VPOS<525)THEN
	   HPOS<=0;
		VPOS<=VPOS+1;
	ELSE
		VPOS<=0;
	END IF;

	IF ((HPOS>656) AND (HPOS<752)) THEN
		HSYNC <='0';
	ELSE
		HSYNC <= '1';
	END IF;
	
	IF ((VPOS>490) AND (VPOS<492)) THEN
		VSYNC <='0';
	ELSE
		VSYNC <= '1';
	END IF;
	
	IF((HPOS>640) OR (VPOS>480))THEN
		R<=(OTHERS=>'0');
		G<=(OTHERS=>'0');
		B<=(OTHERS=>'0');
	END IF;	

END IF;
    

END PROCESS;
END MAIN;


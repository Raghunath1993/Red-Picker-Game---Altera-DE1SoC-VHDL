library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

PACKAGE SCREEN IS
PROCEDURE DISPLAY(SIGNAL XCUR,YCUR:IN INTEGER;
SIGNAL R,G,B:OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END SCREEN;
PACKAGE BODY SCREEN IS
 PROCEDURE DISPLAY(SIGNAL XCUR,YCUR:IN INTEGER;
SIGNAL R,G,B:OUT STD_LOGIC_VECTOR(7 DOWNTO 0)) IS 
BEGIN
IF((XCUR>110 AND XCUR<210) AND(YCUR>70 AND YCUR<170)) THEN
	R<=(OTHERS=>'1');
	G<=(OTHERS=>'1');
	B<=(OTHERS=>'0');
END IF;
IF((XCUR>110 AND XCUR<210) AND(YCUR>310 AND YCUR<410)) THEN
	R<=(OTHERS=>'1');
	G<=(OTHERS=>'0');
	B<=(OTHERS=>'0');
END IF;
IF((XCUR>430 AND XCUR<530) AND(YCUR>70 AND YCUR<170)) THEN
	R<=(OTHERS=>'1');
	G<=(OTHERS=>'1');
	B<=(OTHERS=>'1');
END IF;
IF((XCUR>430 AND XCUR<530) AND(YCUR>310 AND YCUR<410)) THEN
	R<=(OTHERS=>'1');
	G<=(OTHERS=>'0');
	B<=(OTHERS=>'1');
END IF;
END DISPLAY;
END SCREEN;